module divison(
    input        clk,
    input [31:0] src1, rsc2;

);

	// ------------------------------ Division ------------------------------- //
	reg [31:0] dividend;
	reg [62:0] divisor;
	reg [31:0] quotient, quotient_msk;

	reg div_sign;
	reg div_busy = 1'b0;
	reg div_finished = 1'b0;

	wire 


endmodule