// Nosso processador 
module franken_riscv(
			  input  		     clk, reset,
           output reg [31:0] pc,
           input      [31:0] instruction,
           output 		     mem_write,
			  output     [3: 0] byte_enable,
           output     [31:0] alu_result, 
			  output     [31:0] write_data,
           input      [31:0] read_data
	);

	// Registradores
	wire [31:0] src1;
	wire [31:0] src2;
	wire [31:0] data_load;

	//JUMP
	wire is_conditional_jump;
	wire [31:0] jump_add;

	//PC
	wire [31:0] next_pc;
	
	// Atualiza nosso valor de PC
	assign next_pc =	reset 					? 32'b0:
							is_conditional_jump	? jump_add:
							pc + 32'd4;
						  
	always @(posedge clk)
     pc <= next_pc;
	
	// Recebe os valores que sao passados na instruçao
	wire [6:0] opcode;
	assign opcode = instruction[6:0];
	wire [4:0] rd_;
	assign rd_ = instruction[11:7];
	wire [2:0] funct3_;
	assign funct3_ = instruction[14:12];
	wire [4:0] rs1;
	assign rs1 = instruction[19:15];
	wire [4:0] rs2;
	assign rs2 = instruction[24:20];
	wire [6:0] funct7_;
	assign funct7_ = instruction[31:25];
	
	//Instruction Type 
	wire R_type;
	assign R_type = (opcode == 7'b0110011);
	
	wire I_type;
	assign I_type = (opcode == 7'b1100111 | opcode == 7'b0000011 | opcode == 7'b0010011); //Tambem seria uma instruçao do tipo I para 64bits => 0010011
	
	wire S_type;
	assign S_type = (opcode == 7'b0100011); //Tambem seria uma instruçao do tipo S para Double ou Float => 0100111
	
	wire B_type;
	assign B_type = (opcode == 7'b1100011);
	
	wire U_type;
	assign U_type = (opcode == 7'b0110111 | opcode == 7'b0010111);
	
	wire J_type;
	assign J_type = (opcode == 7'b1101111);
	
	// Decodificaçao das instruçoes e seus respectivos tipos 
	wire [4:0] RS1;
	assign RS1 = (R_type | I_type | S_type | B_type) 	? rs1 : 5'b0;
	
	wire [4:0] RS2;
	assign RS2 = (R_type | S_type | B_type)         	? rs2 : 5'b0;

	wire [4:0] RD;
	assign RD = (R_type | I_type | U_type | J_type) 	? rd_ : 5'b0;
	
	wire [2:0] funct3;
	assign funct3 = (R_type | I_type | S_type | B_type)? funct3_ : 3'b0;
	
	wire [6:0] funct7;
	assign funct7 = (R_type)                           ? funct7_ : 7'b0;
	
	wire [31:0] imm;
	assign imm = (I_type) ? ({{20{instruction[31]}},instruction[31:20]}):
					 (S_type) ? ({{20{instruction[31]}},instruction[31:25],instruction[11:7]}):		
					 (B_type) ? ({{19{instruction[31]}},instruction[31],instruction[7],instruction[30:25],instruction[11:8],1'b0}):
					 (U_type) ? ({instruction[31:12],12'b0}):
					 (J_type) ? ({{11{instruction[31]}}, instruction[31],instruction[19:12],instruction[20],instruction[30:21],1'b0}):
					 32'b0;
					 
	//Math
	wire is_add;
	assign is_add    	= (opcode == 7'b0110011 & funct3 == 3'b000 & funct7 == 7'b0000000);
	
	wire is_addi;
	assign is_addi   	= (opcode == 7'b0010011 & funct3 == 3'b000);
	
	wire is_sub;
	assign is_sub 	  	= (opcode == 7'b0110011 & funct3 == 3'b000 & funct7 == 7'b0100000);
	
	//Logic
	wire is_xor;
	assign is_xor	 	= (opcode == 7'b0110011 & funct3 == 3'b100 & funct7 == 7'b0000000);
	
	wire is_or;
	assign is_or	 	= (opcode == 7'b0110011 & funct3 == 3'b110 & funct7 == 7'b0000000);
	
	wire is_andi;
	assign is_andi		= (opcode == 7'b0010011 & funct3 == 3'b111);
	
	//Bit operator
	wire is_slli;
	assign is_slli   	= (opcode == 7'b0010011 & funct3 == 3'b001 & funct7 == 7'b0000000);
	
	wire is_srli;
	assign is_srli	 	= (opcode == 7'b0010011 & funct3 == 3'b101 & funct7 == 7'b0000000);
	
	//PC operator 
	wire is_auipc;
	assign is_auipc  	= (opcode == 7'b0010111);
	
	//Jump 
	wire is_jal;
	assign is_jal    	= (opcode == 7'b1101111);
	
	wire is_lui;
	assign is_lui	  	= (opcode == 7'b0110111);
	
	wire is_jalr;
	assign is_jalr   	= (opcode == 7'b1100111 & funct3 == 3'b0);
	
	wire is_bge;
	assign is_bge    	= (opcode == 7'b1100011 & funct3 == 3'b101);
	
	wire is_beq;
	assign is_beq    	= (opcode == 7'b1100011 & funct3 == 3'b0);
	
	wire is_blt;
	assign is_blt    	= (opcode == 7'b1100011 & funct3 == 3'b100);
	
	wire is_bne;
	assign is_bne    	= (opcode == 7'b1100011 & funct3 == 3'b001);
	
	//Memory 
	wire is_sw;
	assign is_sw     	= (opcode == 7'b0100011 & funct3 == 3'b010);
	
	wire is_lw;
	assign is_lw     	= (opcode == 7'b0000011 & funct3 == 3'b010);
	
	wire is_sb;
	assign is_sb		= (opcode == 7'b0100011 & funct3 == 3'b000);
	
	wire is_lbu;
	assign is_lbu		= (opcode == 7'b0000011 & funct3 == 3'b100);

	//---------------------------- Controler ---------------------------------------------//
	
	parameter   FETCH   = 4'b0000; 	// State 0
   parameter   DECODE  = 4'b0001; 	// State 1
   parameter   MEMADR  = 4'b0010;	// State 2
   parameter   MEMRD   = 4'b0011;	// State 3
   parameter   MEMWB   = 4'b0100;	// State 4
   parameter   MEMWR   = 4'b0101;	// State 5
   parameter   RTYPEEX = 4'b0110;	// State 6
   parameter   ITYPEEX = 4'b0111;	// State 7
   parameter   JEX     = 4'b1000;	// State 8
   parameter   ALUWB   = 4'b1001;	// State 9
   parameter   BEQX    = 4'b1010;	// state 10
	
	wire is_mem_reg;
	wire reg_write;
	wire [3:0] current_state;
	reg  [3:0] next_state;
	
	always @(posedge clk)
		if(reset) current_state <= FETCH;
		else current_state <= next_state;
	
	//Condiçao de escrita na memoria
	assign mem_write = S_type;
	
	//Condiçao de salto
	assign is_conditional_jump = (is_beq || is_bne || is_blt || is_bge || is_jal || is_jalr);
	
	//Escrita da memoria para o registrador
	assign is_mem_reg = is_lw || is_lbu;
	
	// Condicional para escrita nos registradores
	assign reg_write = (R_type || S_type || B_type || I_type || U_type) && RD != 5'b0;
	
	always @*
	begin
		case(current_state)
			FETCH: next_state <= DECODE;
			DECODE: next_state <= (S_type) ? MEMADR : 
                               (R_type) ? RTYPEEX:
										 (I_type) ? ITYPEEX:
										 (J_type) ? JEX:
										 (is_beq || bge || blt
	
	
	end
	
	
	//-------------------------------------ALU-------------------------------------------------//
	wire [31:0] result;
	assign result = 	is_add   	? src1 + src2:
							is_addi		? src1 + imm:
							is_sub		? src1 - src2:
							is_andi		? src1 & imm:
							is_or			? src1 | src2:
							is_slli		? src1 << imm[4:0]:
							is_srli		? src1 >> imm[4:0]:
							is_auipc		? pc + $signed(imm):
							J_type   	? jump_add:
							S_type 		? src1 + imm: 
							is_lw			? src1 + imm: 
							is_sw			? src1 + imm: 
							is_lui		? imm:
							is_xor		? src1 ^ src2:
							is_lbu		? src1 + imm:
							32'b0;
							
	// Recebe o resultado da alu.
	assign alu_result = result;
	
	// Caso nossa instruçao seja de JUMP, temos que calcular a nova posiçao para nosso PC.
	assign jump_add =	is_jal  													? pc 					+ $signed(imm):
							is_jalr 													? $signed(src1) 	+ $signed(imm):
							(is_beq && ($signed(src1) == $signed(src2))) ? pc		 			+ $signed(imm) :
							(is_bne && ($signed(src1) != $signed(src2))) ? pc 					+ $signed(imm):
							(is_blt && ($signed(src1)  < $signed(src2)))	? pc			 		+ $signed(imm):
							(is_bge && ($signed(src1) >= $signed(src2)))	? pc 					+ $signed(imm):
							pc + 32'd4;

	// Valor que sera salvo na nossa memoria e a condicional de escrita
	assign write_data = is_sw ? src2 : (is_sb ? (alu_result[1:0]==3 ? {src2[7:0], 24'h000000} : 
														      alu_result[1:0]==2 ? {8'h00, src2[7:0], 16'h0000} :
														      alu_result[1:0]==1 ? {16'h0000, src2[7:0], 8'h00} :
														                           {24'h000000, src2[7:0]}) :
																							32'bX);
	
	// Escrita alinhada na memoria
	assign byte_enable = is_lbu || is_sb ? (alu_result[1:0]==3 ? 4'b1000 : // sb/lb
														 alu_result[1:0]==2 ? 4'b0100 :
														 alu_result[1:0]==1 ? 4'b0010 :
														                      4'b0001): 
														                      4'b1111;  // lw/sw
	
   //Acerta a posiçao para ser salvo em memoria 
   assign data_load = is_lbu ? (alu_result[1:0]==3 ? {24'h000000, read_data[31:24]} : 
	                             alu_result[1:0]==2 ? {24'h000000, read_data[23:16]} : 
	                             alu_result[1:0]==1 ? {24'h000000, read_data[15: 8]} : 
										                       {24'h000000, read_data[ 7: 0]}):
																	  read_data;
	
	regfile regs(clk, reg_write, RS1, RS2, RD, is_mem_reg ? data_load : alu_result, src1, src2);
	
endmodule

module control_unit(input wire       clk,
						  input wire [6:0] opcode,
						  input wire [2:0] funct3,
						  input wire [6:0] funct7);
						  
						  

endmodule

// Modulo de registradores
module regfile(input  wire        clk, 
               input  wire        reg_write,
               input  wire [4:0]  reg_addr1, reg_addr2, addr, 
               input  wire [31:0] write_reg, 
               output wire [31:0] rd1, rd2);
					
  reg [31:0] rf[31:0];

	always @(posedge clk) 
		if (reg_write) 
			rf[addr] <= write_reg;	
		
	assign rd1 = (reg_addr1 != 32'b0) ? rf[reg_addr1] : 32'b0; 
	assign rd2 = (reg_addr2 != 32'b0) ? rf[reg_addr2] : 32'b0;
endmodule